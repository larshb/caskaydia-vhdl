--  ===>
--  ==>
--  =>
--  <=
--  <==
--  <===
